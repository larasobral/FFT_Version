module memory_ed2 #(parameter W = 16, parameter N = 16)(
	output reg signed [7:0] sin_rom[16:0],
	output reg signed [7:0] cos_rom[16:0]);

	initial 
	   begin 

		sin_rom[0] = 17'b0_0000000000000000;
		cos_rom[0] = 17'b0_1000000000000000;

		sin_rom[1] = 17'b0_0011101100111100;  
		cos_rom[1] = 17'b0_1110110011110010; 

		sin_rom[2] = 17'b0_0111100000000000; 
		cos_rom[2] = 17'b0_1000000000000000; 

		sin_rom[3] = 17'b0_1011010101011011; 
		cos_rom[3] = 17'b0_0110101010101101; 

		sin_rom[4] = 17'b0_1100000000000000;  
		cos_rom[4] = 17'b0_0000000000000000;  
 
		sin_rom[5] = 17'b0_1011010101011011;   
		cos_rom[5] = 17'b0_1001010101011011;  

		sin_rom[6] = 17'b0_0111100000000000;  
		cos_rom[6] = 17'b0_0111111111111111;  
 
		sin_rom[7] = 17'b0_0011101100111100;   
		cos_rom[7] = 17'b0_1011011000111000; 

		sin_rom[8] = 17'b1_0000000000000000; 
		cos_rom[8] = 17'b1_1000000000000000; 

		sin_rom[9] = 17'b1_0101101100111100;  
		cos_rom[9] = 17'b1_0101100111100111;  

		sin_rom[10] = 17'b1_1000000000000000; 
		cos_rom[10] = 17'b1_0000000000000000;  

		sin_rom[11] = 17'b1_1101100111100000;  
		cos_rom[11] = 17'b1_1001100111100111; 

		sin_rom[12] = 17'b1_1110000000000000;  
		cos_rom[12] = 17'b1_0111111111111111;  

		sin_rom[13] = 17'b1_1101100111100000; 
		cos_rom[13] = 17'b1_0011010101011010;  

		sin_rom[14] = 17'b1_1011010101011011; 
		cos_rom[14] = 17'b1_0000000000000000;  

		sin_rom[15] = 17'b1_1000000000000000; 
		cos_rom[15] = 17'b1_1001011000111000; 

		sin_rom[16] = 17'b1_0111100000000000;  
		cos_rom[16] = 17'b1_1000000000000000;  

		sin_rom[17] = 17'b1_0000000000000000;  
		cos_rom[17] = 17'b1_0111111111111111; 

		sin_rom[20] = 17'b1_1100000000000000;   
		cos_rom[20] = 17'b1_0000000000000000; 

		sin_rom[21] = 17'b1_1011010101011011;    
		cos_rom[21] = 17'b1_0101101010101100;  

		sin_rom[22] = 17'b1_0111100000000000;   
		cos_rom[22] = 17'b1_1000000000000000; 

		sin_rom[24] = 17'b0_0000000000000000;    
		cos_rom[24] = 17'b1_1100000000000000; 

		sin_rom[25] = 17'b0_0011101100111100;  
		cos_rom[25] = 17'b1_0011100111100111; 

		sin_rom[26] = 17'b0_0101101100111100;  
		cos_rom[26] = 17'b1_1010101010101100; 

		sin_rom[27] = 17'b0_0111000000000000;  
		cos_rom[27] = 17'b1_0111000000000000; 
  
		sin_rom[28] = 17'b0_0110000000000000;  
		cos_rom[28] = 17'b1_0000000000000000; 

		sin_rom[30] = 17'b0_0101000000000000;  
		cos_rom[30] = 17'b1_1000000000000000;  

		sin_rom[32] = 17'b0_0100000000000000;  
		cos_rom[32] = 17'b1_1000000000000000;  

		sin_rom[33] = 17'b0_0010101010101101;   
		cos_rom[33] = 17'b1_0101000000000000;  

		sin_rom[35] = 17'b0_0000100111100111;
		cos_rom[35] = 17'b1_0010101010101011;  

		sin_rom[36] = 17'b0_0000000001111000;  
		cos_rom[36] = 17'b1_0000100111100110; 

		sin_rom[39] = 17'b0_0000000000000000; 
		cos_rom[39] = 17'b1_1111111111111111;  

		sin_rom[40] = 17'b0_0000000000000000; 
		cos_rom[40] = 17'b1_1011010101011010; 

		sin_rom[42] = 17'b0_0000000001111000; 
		cos_rom[42] = 17'b1_0111111111111111;  

		sin_rom[44] = 17'b0_0000100111100111;
		cos_rom[44] = 17'b1_0000000000000000; 

		sin_rom[45] = 17'b0_0000101010101101; 
		cos_rom[45] = 17'b1_1000000001111000;

		sin_rom[48] = 17'b0_0000000000000000;  
		cos_rom[48] = 17'b1_1000000000000000;  

		sin_rom[50] = 17'b0_0000100000000000;   
		cos_rom[50] = 17'b1_0000000001111000;  

		sin_rom[52] = 17'b0_0000101010101101;   
		cos_rom[52] = 17'b1_0101010101011010;  

		sin_rom[54] = 17'b0_0000000001111000; 
		cos_rom[54] = 17'b1_1100000000000000; 

		sin_rom[55] = 17'b0_1000000000001100;  
		cos_rom[55] = 17'b1_0011101100111000; 

		sin_rom[56] = 17'b0_1000000000000000;      
		cos_rom[56] = 17'b1_1000000000000000;  

		sin_rom[60] = 17'b0_1000000000000000;      
		cos_rom[60] = 17'b1_0111111111111111; 

		sin_rom[63] = 17'b0_1000000000001100; 
		cos_rom[63] = 17'b1_1001100111100110; 

		sin_rom[64] = 17'b0_1000000000000000; 
		cos_rom[64] = 17'b1_0110101010101011;  

		sin_rom[65] = 17'b0_1000000000001100;  
		cos_rom[65] = 17'b1_1001011000110110;  

		sin_rom[66] = 17'b0_1000000000000000;    
		cos_rom[66] = 17'b1_1000000000000000; 

		sin_rom[70] = 17'b0_1000000000000000;       
		cos_rom[70] = 17'b1_0000000000000000; 

		sin_rom[72] = 17'b0_1000000000000000;  
		cos_rom[72] = 17'b1_0000000000000000;  

		sin_rom[75] = 17'b0_1000000000001100;   
		cos_rom[75] = 17'b1_0000000000000000; 

		sin_rom[77] = 17'b0_1000000000000000;     
		cos_rom[77] = 17'b1_0000000000000000;  

		sin_rom[78] = 17'b0_1000000000000000; 
		cos_rom[78] = 17'b1_0000000000000000;  

		sin_rom[80] = 17'b0_1000000000000000;  
		cos_rom[80] = 17'b1_1011010101011001; 

		sin_rom[81] = 17'b0_1000000000000000;
		cos_rom[81] = 17'b1_1000000001111000;  

		sin_rom[84] = 17'b0_1000000000001100; 
		cos_rom[84] = 17'b1_0111111111111111; 

		sin_rom[88] = 17'b0_1000000000000000; 
		cos_rom[88] = 17'b1_0000000111011111;  

		sin_rom[90] = 17'b0_1000000000000000;  
		cos_rom[90] = 17'b1_1000000000001101; 

		sin_rom[91] = 17'b0_1000000000001100; 
		cos_rom[91] = 17'b1_1000000000000000; 

		sin_rom[96] = 17'b0_1000000000000000; 
		cos_rom[96] = 17'b1_1000000000000000; 

		sin_rom[98] = 17'b0_1000000000001100; 
		cos_rom[98] = 17'b1_1000000000000000; 

		sin_rom[99] = 17'b0_1000000000000000;  
		cos_rom[99] = 17'b1_1000000000000000;  

		sin_rom[100] = 17'b0_1000000000000000;    
		cos_rom[100] = 17'b1_1000000000000000;  

		sin_rom[104] = 17'b0_1000000000000000;   
		cos_rom[104] = 17'b1_1000000000001101; 

		sin_rom[105] = 17'b0_1000000000000000; 
		cos_rom[105] = 17'b1_1000000000001101;

		sin_rom[108] = 17'b0_1000000000001100;    
		cos_rom[108] = 17'b1_1000000000000000;

		sin_rom[110] = 17'b0_1000000000000000;  
		cos_rom[110] = 17'b1_1000000000000000;
         
		sin_rom[112] = 17'b0_1000000000000000;   
		cos_rom[112] = 17'b1_1000000000000000;

		sin_rom[117] = 17'b0_1000000000000000;      
		cos_rom[117] = 17'b1_1000000000000000;

		sin_rom[120] = 17'b0_1000000000001100; 
		cos_rom[120] = 17'b1_1000000001111000;  

		sin_rom[121] = 17'b0_1000000000000000;  
		cos_rom[121] = 17'b1_1000000011011000;  

		sin_rom[126] = 17'b0_1000000000000000; 
		cos_rom[126] = 17'b1_1000000000000000; 

		sin_rom[130] = 17'b0_1000000000000000;  
		cos_rom[130] = 17'b1_1000000000000000; 

		sin_rom[132] = 17'b0_1000000000000000;
		cos_rom[132] = 17'b1_1000000000000000;  

		sin_rom[135] = 17'b0_1000000000000000;  
		cos_rom[135] = 17'b1_1000000000000000; 

		sin_rom[140] = 17'b0_1000000000001100;  
		cos_rom[140] = 17'b1_1000000000000000;  

		sin_rom[143] = 17'b0_1000000000000000;    
		cos_rom[143] = 17'b1_1000000000000000; 

		sin_rom[144] = 17'b0_1000000000000000;
		cos_rom[144] = 17'b1_1000000000000000;  

		sin_rom[150] = 17'b0_1000000000000000;    
		cos_rom[150] = 17'b1_1000000000000000; 

		sin_rom[154] = 17'b0_1000000000001100;     
		cos_rom[154] = 17'b1_1000000000000000; 

		sin_rom[156] = 17'b0_1000000000000000;   
		cos_rom[156] = 17'b1_1000000000000000; 

		sin_rom[165] = 17'b0_1000000000000000;    
		cos_rom[165] = 17'b1_1000000000000000; 

		sin_rom[168] = 17'b0_1000000000000000;   
		cos_rom[168] = 17'b1_1000000000000000; 

		sin_rom[169] = 17'b0_1000000000001100;   
		cos_rom[169] = 17'b1_1000000000000000;

		sin_rom[180] = 17'b0_1000000000000000; 
		cos_rom[180] = 17'b1_1000000000000000;

		sin_rom[182] = 17'b0_1000000000000000; 
		cos_rom[182] = 17'b1_1000000000000000; 

		sin_rom[195] = 17'b0_1000000000001100;   
		cos_rom[195] = 17'b1_1000000000001111;

		sin_rom[196] = 17'b0_1000000000000000;  
		cos_rom[196] = 17'b1_1000000000001111;

		sin_rom[210] = 17'b0_1000000000000000; 
		cos_rom[210] = 17'b1_1000000000000000;

		sin_rom[225] = 17'b0_1000000000001100; 
		cos_rom[225] = 17'b1_1000000001111000;
           end

endmodule
